module def();
    `define HOLD 2'b00
    `define RESET 2'b01
    `define SET 2'b10
    `define TOGGLE 2'b11
endmodule