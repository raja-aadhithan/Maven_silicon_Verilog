module fifo_tb();
reg clk,aresetn,read,write;
reg [7:0]data_in;
wire full,empty;
wire [7:0]data_out;
integer i;

fifo dut(clk,aresetn,read,write,data_in,full,empty,data_out);
initial begin 
    clk = 1'b1;
    forever #5 clk = ~clk;
end

initial begin
    $monitor("$@time:%3d, read :%b, write :%b, datain = %b, dataout = %b",$time,read,write,data_in,data_out);
    aresetn = 0;
    #20;
    aresetn = 1;
    write = 1;
    read = 0;
    data_in = 8'd5;
    #10;
    data_in = 8'd15;
    #10;
    data_in = 8'd21;
    #10;
    data_in = 8'd31;
    #10;
    data_in = 8'd41;
    #10;
    data_in = 8'd12;
    #10;
    data_in = 8'd13;
    #10;
    data_in = 8'd33;
    #10;
    data_in = 8'd42;
    #10;
    data_in = 8'd16;
    #10;
    read = 1;
    data_in = 8'd2;
    #10;
    data_in = 8'd1;
    #10;
    data_in = 8'd2;
    #10;
    data_in = 8'd3;
    #10;
    data_in = 8'd4;
    #10;
    data_in = 8'd21;
    #10;
    data_in = 8'd31;
    #10;
    data_in = 8'd41;
    #10;
    data_in = 8'd12;
    #10;
    data_in = 8'd13;
    #10;
    data_in = 8'd21;
    #10;
    data_in = 8'd31;
    #10;
    data_in = 8'd41;
    #10;
    data_in = 8'd12;
    #10;
    data_in = 8'd13;
    #10;
    write = 0;
    #30;
    read = 0;
    write =1;
    data_in = 8'd10;
    #10;
    data_in = 8'd11;
    #10;
    data_in = 8'd21;
    #10;
    data_in = 8'd31;
    #10;
    data_in = 8'd41;
    #10;
    data_in = 8'd12;
    #10;
    data_in = 8'd13;
    #10;
    data_in = 8'd33;
    #10;
    data_in = 8'd42;
    #10;
    data_in = 8'd16;
    #10;
    data_in = 8'd22;
    #10;
    data_in = 8'd30;
    #10;
    data_in = 8'd06;
    #10;
    read = 1;
    write = 0;
    #35;
    write =1;
    data_in = 8'd30;
    #10;
    data_in = 8'd06;
    write =0;
    #500;
    $finish;
end
endmodule